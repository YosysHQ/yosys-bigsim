@0000000  98 00 00 00 78 1c 00 00 3b 9c ff fc b8 00 d8 00
@0000010  78 01 00 00 38 21 81 80 78 02 00 00 38 42 81 88
@0000020  4c 22 00 04 58 20 00 00 34 21 00 04 e3 ff ff fd
@0000030  f8 00 00 53 78 01 de ad 38 02 be ef 58 22 00 00
@0000040  37 9c ff e8 5b 8b 00 14 5b 8c 00 10 5b 8d 00 0c
@0000050  5b 9b 00 08 5b 9d 00 04 34 1b 00 18 b7 7c d8 00
@0000060  5b 61 00 00 2b 61 00 00 34 02 00 05 f8 00 00 a5
@0000070  b8 20 68 00 78 0b 00 00 39 6b 81 80 34 02 00 02
@0000080  f8 00 00 78 b5 61 08 00 28 2b 00 00 2b 61 00 00
@0000090  20 22 00 1f 34 01 00 01 f8 00 00 72 b9 61 60 00
@00000a0  78 0b 00 00 39 6b 81 80 b9 a0 08 00 34 02 00 02
@00000b0  f8 00 00 6c b5 61 08 00 58 2c 00 00 2b 8b 00 14
@00000c0  2b 8c 00 10 2b 8d 00 0c 2b 9b 00 08 2b 9d 00 04
@00000d0  37 9c 00 18 c3 a0 00 00 37 9c ff f0 5b 8b 00 0c
@00000e0  5b 9b 00 08 5b 9d 00 04 34 1b 00 10 b7 7c d8 00
@00000f0  5b 61 00 00 2b 61 00 00 34 02 00 05 f8 00 00 81
@0000100  78 0b 00 00 39 6b 81 80 34 02 00 02 f8 00 00 55
@0000110  b5 61 08 00 28 2b 00 00 2b 61 00 00 20 22 00 1f
@0000120  34 01 00 01 f8 00 00 4f a1 61 08 00 7c 21 00 00
@0000130  2b 8b 00 0c 2b 9b 00 08 2b 9d 00 04 37 9c 00 10
@0000140  c3 a0 00 00 37 9c ff f4 5b 9b 00 08 5b 9d 00 04
@0000150  34 1b 00 0c b7 7c d8 00 5b 61 00 00 78 01 ff 00
@0000160  38 21 00 04 2b 62 00 00 58 22 00 00 2b 9b 00 08
@0000170  2b 9d 00 04 37 9c 00 0c c3 a0 00 00 37 9c ff ec
@0000180  5b 9b 00 08 5b 9d 00 04 34 1b 00 14 b7 7c d8 00
@0000190  34 01 00 02 fb ff ff ec 34 01 00 00 5b 61 ff f8
@00001a0  e0 00 00 28 2b 61 ff f8 fb ff ff cc b8 20 10 00
@00001b0  34 01 00 00 5c 41 00 20 2b 61 ff f8 b4 21 08 00
@00001c0  34 21 00 03 fb ff ff e0 2b 61 ff f8 34 02 00 02
@00001d0  f8 00 00 24 34 21 00 06 5b 61 ff fc 2b 61 ff fc
@00001e0  20 22 00 01 34 01 00 00 44 41 00 0b 2b 61 ff fc
@00001f0  34 21 ff fd 34 02 00 01 f8 00 00 42 5b 61 00 00
@0000200  2b 62 00 00 34 01 00 3f 54 41 00 0b 2b 61 00 00
@0000210  fb ff ff 8c 2b 61 ff f8 b4 21 08 00 b8 20 10 00
@0000220  2b 61 ff fc b4 41 08 00 34 21 00 03 5b 61 ff fc
@0000230  e3 ff ff eb 2b 61 ff f8 34 21 00 01 5b 61 ff f8
@0000240  2b 62 ff f8 34 01 00 3f 50 22 ff d7 34 01 00 00
@0000250  2b 9b 00 08 2b 9d 00 04 37 9c 00 14 c3 a0 00 00
@0000260  20 42 00 1f 78 03 00 00 38 63 80 00 b4 42 10 00
@0000270  b4 42 10 00 b4 62 18 00 28 63 00 00 c0 60 00 00
@0000280  b4 21 08 00 b4 21 08 00 b4 21 08 00 b4 21 08 00
@00002f0  b4 21 08 00 b4 21 08 00 b4 21 08 00 c3 a0 00 00
@0000300  20 42 00 1f 78 03 00 00 38 63 80 80 b4 42 10 00
@0000310  b4 42 10 00 b4 62 18 00 28 63 00 00 c0 60 00 00
@0000320  00 21 00 01 00 21 00 01 00 21 00 01 00 21 00 01
@0000390  00 21 00 01 00 21 00 01 00 21 00 01 c3 a0 00 00
@00003a0  20 42 00 1f 78 03 00 00 38 63 81 00 b4 42 10 00
@00003b0  b4 42 10 00 b4 62 18 00 28 63 00 00 c0 60 00 00
@00003c0  14 21 00 01 14 21 00 01 14 21 00 01 14 21 00 01
@0000430  14 21 00 01 14 21 00 01 14 21 00 01 c3 a0 00 00
@0000440  00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
@0008000  00 00 02 fc 00 00 02 f8 00 00 02 f4 00 00 02 f0
@0008010  00 00 02 ec 00 00 02 e8 00 00 02 e4 00 00 02 e0
@0008020  00 00 02 dc 00 00 02 d8 00 00 02 d4 00 00 02 d0
@0008030  00 00 02 cc 00 00 02 c8 00 00 02 c4 00 00 02 c0
@0008040  00 00 02 bc 00 00 02 b8 00 00 02 b4 00 00 02 b0
@0008050  00 00 02 ac 00 00 02 a8 00 00 02 a4 00 00 02 a0
@0008060  00 00 02 9c 00 00 02 98 00 00 02 94 00 00 02 90
@0008070  00 00 02 8c 00 00 02 88 00 00 02 84 00 00 02 80
@0008080  00 00 03 9c 00 00 03 98 00 00 03 94 00 00 03 90
@0008090  00 00 03 8c 00 00 03 88 00 00 03 84 00 00 03 80
@00080a0  00 00 03 7c 00 00 03 78 00 00 03 74 00 00 03 70
@00080b0  00 00 03 6c 00 00 03 68 00 00 03 64 00 00 03 60
@00080c0  00 00 03 5c 00 00 03 58 00 00 03 54 00 00 03 50
@00080d0  00 00 03 4c 00 00 03 48 00 00 03 44 00 00 03 40
@00080e0  00 00 03 3c 00 00 03 38 00 00 03 34 00 00 03 30
@00080f0  00 00 03 2c 00 00 03 28 00 00 03 24 00 00 03 20
@0008100  00 00 04 3c 00 00 04 38 00 00 04 34 00 00 04 30
@0008110  00 00 04 2c 00 00 04 28 00 00 04 24 00 00 04 20
@0008120  00 00 04 1c 00 00 04 18 00 00 04 14 00 00 04 10
@0008130  00 00 04 0c 00 00 04 08 00 00 04 04 00 00 04 00
@0008140  00 00 03 fc 00 00 03 f8 00 00 03 f4 00 00 03 f0
@0008150  00 00 03 ec 00 00 03 e8 00 00 03 e4 00 00 03 e0
@0008160  00 00 03 dc 00 00 03 d8 00 00 03 d4 00 00 03 d0
@0008170  00 00 03 cc 00 00 03 c8 00 00 03 c4 00 00 03 c0
